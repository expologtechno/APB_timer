`include "base_seq.sv"
`include "reset_seq.sv"
`include "sanity_seq.sv"

`include "base_seq.sv"

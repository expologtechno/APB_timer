//======================= TRANSACTION =====================================/
class output_transaction extends uvm_sequence_item;

`uvm_object_utils(output_transaction)


      
//--------------------------constructor--------------------------------	
function new(string name="output_transaction");
super.new(name);
endfunction


endclass

`include "interface.sv"

`include "../agent/apb_agent/apb_transaction.sv"
`include "../agent/apb_agent/apb_driver.sv"
`include "../agent/apb_agent/apb_monitor.sv"
`include "../agent/apb_agent/apb_sequencer.sv"
`include "../agent/apb_agent/apb_agent.sv"


`include "../agent/reset_agent/reset_tx.sv"
`include "../agent/reset_agent/reset_driver.sv"
`include "../agent/reset_agent/reset_sequencer.sv"
`include "../agent/reset_agent/reset_agent.sv"

`include "../agent/passive_agent/output_tx.sv"
`include "../agent/passive_agent/output_monitor.sv"
`include "../agent/passive_agent/output_agent.sv"


`include "virtual_sequencer.sv"
`include "../seqs/seq_list.svh"

`include "virtual_sequence.sv"

`include "scoreboard.sv"
`include "env.sv"

`include "../test/test_list.svh"

`include "base_test.sv"

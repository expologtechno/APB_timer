`include "base_test.sv"
`include "reset_test.sv"
`include "sanity_test.sv"
